// This file declares all uvm libs and uvm macros

`ifndef PACK_SV
`define PACK_SV

`include "uvm_macros.svh"
import uvm_pkg::*;

`endif 